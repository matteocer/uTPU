parameter int ARRAY_SIZE = 2;
parameter int INPUT_DATA_WIDTH = 4;
parameter int ACCUMULATOR_DATA_WIDTH = 16;
